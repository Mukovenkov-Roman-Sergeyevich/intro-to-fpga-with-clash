../../../src/05-bus/merge_serial_to_parallel.sv