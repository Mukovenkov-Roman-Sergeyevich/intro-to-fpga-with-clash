../../../src/05-bus/serial_to_parallel/serial_to_parallel.sv