../../../src/05-bus/merge_parallel/merge_parallel.sv